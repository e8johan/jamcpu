-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package p0_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 10;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"00000100001000000000000000111000",
		"00000100010000001111111100100110",
		"11110000011000000000000000000000",
		"00001000001000011111111111111100",
		"00001000010000100000000000000001",
		"01000100011000110000000000001000",
		"10110000100000010000000000000000",
		"01100000101000010001000000000000",
		"01011100101000000000000000000000",
		"00000000000000000000000000000000");
end;