-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package p1_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 25;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"00000000000000000000000000000000",
		"01111111110000000000000000001110",
		"00000100001000000000000000001100",
		"00000000100000000000000000000000",
		"10001100010000010000000100000000",
		"10001100011000010000000100000100",
		"00100000101000100001100000000000",
		"00000100001000011111111111111100",
		"00000000100001000010100000000000",
		"01100000101000000000100000000000",
		"01011100101000001111111111111010",
		"00000000000000000000000000000000",
		"10011100100000000000000100001000",
		"01001100000000000000000000000000",
		"00000000000000000000000000000000",
		"00000100001000000000000000100000",
		"10011100001000010000000011111111",
		"00000100001000011111111111111100",
		"01011100001000001111111111111110",
		"00000000000000000000000000000000",
		"01111100000111100000000000000001",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000");
end;