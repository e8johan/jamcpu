-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package sni_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 58;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"11110001011000000000000000000000",
		"00000101100000001111111100000000",
		"01010001100010110000000000000100",
		"00000000000000000000000000000000",

		"11110100000000001111101100000000",
		"01111100000000000000000000001001",
		"00000101100010111111101100000000",
		"01111100000111110000000000000000",

		"00000100001000000000000000101010",
		"10011100001000000000000000000000",
		"00000100001000000000000000000001",
		"10011100001000000000000000000001",

		"00000100001000000000000000110111",
		"10011100001000000000000000000010",
		"00000100001000000000000000000111",
		"10011100001000000000000000000011",

		"00000100001000000000000000001001",
		"10011100001000000000000000000100",
		"00000100001000000000000000001101",
		"10011100001000000000000000000101",

		"00000100001000000000000000111111",
		"10011100001000000000000000000110",
		"00000100001000000000000000010011",
		"10011100001000000000000000000111",

		"00000100001000000000000000000010",
		"10011100001000000000000000001000",
		"00000100001000000000000000000011",
		"10011100001000000000000000001001",

		"00000100001000000000000000000100",
		"10011100001000000000000000001010",
		"00000100001000000000000001011001",
		"10011100001000000000000000001011",

		"00000100001000000000000000111101",
		"10011100001000000000000000001100",
		"00000100001000000000000000101010",
		"10011100001000000000000000001101",

		"00000100001000000000000000000111",
		"10011100001000000000000000001110",
		"00000100001000000000000000001011",
		"10011100001000000000000000001111",

		"00000100001000000000000000000000",
		"00001100010000010000000000000001",
		"10001100011000010000000000000000",
		"10001100100000100000000000000000",

		"01100000101001000001100000000000",
		"01001100101000000000000000000001",
		"00000000000000000000000000000000",
		"10011100011000100000000000000000",

		"10011100100000010000000000000000",
		"00001100010000100000000000000001",
		"00000100101000000000000001000000",
		"01011100010001011111111111110111",

		"00000000000000000000000000000000",
		"00001100001000010000000000000001",
		"01011100001001011111111111110011",
		"00000000000000000000000000000000",

		"01001100000000000000000000000000",
		"00000000000000000000000000000000");
end;