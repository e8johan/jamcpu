-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package mul_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 10;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"00000000000000000000000000000000",
		"00000100001000000000000000000000",
		"00000100100000000000000000011110",
		"00000100001000010000000000001010",
		"00000100010000010000000000010100",
		"00100000011000100000100000000000",
		"01011100001001001111111111111101",
		"00000100101000000000000000010000",
		"01001100000000000000000000000000",
		"00000000000000000000000000000000");
end;