-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package trap_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 25;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"00000000000000000000000000000000",
		"11100100001000000000000000000000",
		"10110100010000010000001100000000",
		"01001100010000000000000000001101",
		"10110100010000010000001000000000",
		"01100000011000000001000000000000",
		"10001100100000000000000000000000",
		"00000000100001000001100000000000",
		"10011100100000000000000000000000",
		"10110100010000010000000100000000",
		"01100000011000000001000000000000",
		"10001100100000000000000000000001",
		"00000000100001000001100000000000",
		"10011100100000000000000000000000",
		"11110100000000000000001100000000",
		"01111100000111110000000000000001",
		"10011100000000000000000000000000",
		"10011100000000000000000000000001",
		"00000100001000001111111111111111",
		"00001000010000000111111111111111",
		"11000000001000010001000000000000",
		"00010000010000010000100000000000",
		"11111111111111111111111111111111",
		"01001100000000001111111111111011",
		"00000000000000000000000000000000");
end;
