-- ROM package

library ieee;
use ieee.std_logic_1164.all;

package p2_rom is
	constant w:integer:= 32;  --width of ROM
	constant l:integer:= 12;  --lenght of ROM
 	
	subtype rom_word is std_logic_vector(w-1 downto 0);
	type rom_table is array (0 to l-1) of rom_word;

	constant rom_image:rom_table:=rom_table'(
		"11101000001000000000000000000001",
		"00000100010000000000000000000000",
		"00000100011000000000000000000001",
		"00000100100000000000000000010000",
		"10110000101000010001100000000000",
		"01001100101000000000000000001001",
		"00000000000000000000000000000000",
		"10000100110000000001100000000000",
		"01100000101001100000000000000000",
		"01001100101000000000000000000011",
		"00000000000000000000000000000000",
		"00000000110000000000000000000000",
		"10010100110000000010000000000000",
		"01000100011000110000000000000010",
		"01000100100001000000000000000010",
		"00000100010000100000000000000001",
		"01100100101000100000000000000100",
		"01011100101000001111111111110011",
		"00000000000000000000000000000000",
		"11110100000000001000000000000000",
		"01001100000000000000000000000000",
		"00000000000000000000000000000000");
end;